LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY CA2_BCD_8B IS PORT (
	CA2 : IN STD_LOGIC_VECTOR(7 downto 0);
	BCD : OUT STD_LOGIC_VECTOR(7 downto 0));
END CA2_BCD_8B;

ARCHITECTURE taula_veritat OF CA2_BCD_8B IS
	BEGIN	-- nomes hi ha els productes possibles de dos enters entre -56 i 64
	with CA2 SELECT	BCD <= 
		"01100100" WHEN "01000000",  -- 64
		"01010110" WHEN "00111000",  -- 56
		"01001001" WHEN "00110001",  -- 49
		"01001000" WHEN "00110000",  -- 48
		"01000010" WHEN "00101010",  -- 42
		"01000000" WHEN "00101000",  -- 40
		"00110110" WHEN "00100100",  -- 36
		"00110101" WHEN "00100011",  -- 35
		"00110010" WHEN "00100000",  -- 32
		"00110000" WHEN "00011110",  -- 30
		"00101000" WHEN "00011100",  -- 28
		"00100101" WHEN "00011001",  -- 25
		"00100100" WHEN "00011000",  -- 24
		"00100001" WHEN "00010101",  -- 21
		"00100000" WHEN "00010100",  -- 20
		"00011000" WHEN "00010010",  -- 18
		"00010110" WHEN "00010000",  -- 16
		"00010101" WHEN "00001111",  -- 15
		"00010100" WHEN "00001110",  -- 14
		"00010010" WHEN "00001100",  -- 12
		"00010000" WHEN "00001010",  -- 10
		"00001001" WHEN "00001001",  -- 9
		"00001000" WHEN "00001000",  -- 8
		"00000111" WHEN "00000111",  -- 7
		"00000110" WHEN "00000110",  -- 6
		"00000101" WHEN "00000101",  -- 5
		"00000100" WHEN "00000100",  -- 4
		"00000011" WHEN "00000011",  -- 3
		"00000010" WHEN "00000010",  -- 2
		"00000001" WHEN "00000001",  -- 1
		"00000000" WHEN "00000000",  -- 0
		"00000001" WHEN "11111111",  -- -1
		"00000010" WHEN "11111110",  -- -2
		"00000011" WHEN "11111101",  -- -3
		"00000100" WHEN "11111100",  -- -4
		"00000101" WHEN "11111011",  -- -5
		"00000110" WHEN "11111010",  -- -6
		"00000111" WHEN "11111001",  -- -7
		"00001000" WHEN "11111000",  -- -8
		"00001001" WHEN "11110111",  -- -9
		"00010000" WHEN "11110110",  -- -10
		"00010010" WHEN "11110100",  -- -12
		"00010100" WHEN "11110010",  -- -14
		"00010101" WHEN "11110001",  -- -15
		"00010110" WHEN "11110000",  -- -16
		"00011000" WHEN "11101110",  -- -18
		"00100000" WHEN "11101100",  -- -20
		"00100001" WHEN "11101011",  -- -21
		"00100100" WHEN "11101000",  -- -24
		"00100101" WHEN "11100111",  -- -25
		"00101000" WHEN "11100100",  -- -28
		"00110000" WHEN "11100010",  -- -30
		"00110010" WHEN "11100000",  -- -32
		"00110101" WHEN "11011101",  -- -35
		"00110110" WHEN "11011100",  -- -36
		"01000000" WHEN "11011000",  -- -40
		"01000010" WHEN "11010110",  -- -42
		"01001000" WHEN "11010000",  -- -48
		"01001001" WHEN "11001111",  -- -49
		"01010110" WHEN "11001000",  -- -56
		"--------" WHEN OTHERS;
	END taula_veritat;
